
`ifndef __SOC_DEFS__
`define __SOC_DEFS__

`define USE_PLL
`define OUT_IO 8
`define IN_IO 8
`define SSD_OUTPUT
`define NPU_ACCELERATOR

`endif