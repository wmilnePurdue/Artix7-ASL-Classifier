
`ifndef __SOC_DEFS__
`define __SOC_DEFS__

`define USE_PLL
`define GPIO_COUNT 10
//`define SPI_OUTPUT
`define SSD_OUTPUT
`define NPU_ACCELERATOR

`endif